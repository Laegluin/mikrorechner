-- MEM/WB Pipeline Stage

-- entity pipe_mem_wb.vhd

-- WIP
